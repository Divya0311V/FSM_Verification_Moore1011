package fsm_sgls;
 `include "FSM_clk.svh"
 `include "FSM_rst.svh"
 `include "FSM_1.svh"
 `include "FSM_2.svh"
 `include "FSM_3.svh"
 `include "FSM_simulus.svh"
 `include "FSM_runfile.svh"
endpackage
